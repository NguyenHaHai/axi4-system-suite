library verilog;
use verilog.vl_types.all;
entity serv_state is
    generic(
        RESET_STRATEGY  : string  := "MINI";
        WITH_CSR        : vl_logic_vector(0 downto 0) := (others => Hi1);
        ALIGN           : vl_logic_vector(0 downto 0) := (others => Hi0);
        MDU             : vl_logic_vector(0 downto 0) := (others => Hi0);
        W               : integer := 1
    );
    port(
        i_clk           : in     vl_logic;
        i_rst           : in     vl_logic;
        i_new_irq       : in     vl_logic;
        i_alu_cmp       : in     vl_logic;
        o_init          : out    vl_logic;
        o_cnt_en        : out    vl_logic;
        o_cnt0to3       : out    vl_logic;
        o_cnt12to31     : out    vl_logic;
        o_cnt0          : out    vl_logic;
        o_cnt1          : out    vl_logic;
        o_cnt2          : out    vl_logic;
        o_cnt3          : out    vl_logic;
        o_cnt7          : out    vl_logic;
        o_cnt11         : out    vl_logic;
        o_cnt12         : out    vl_logic;
        o_cnt_done      : out    vl_logic;
        o_bufreg_en     : out    vl_logic;
        o_ctrl_pc_en    : out    vl_logic;
        o_ctrl_jump     : out    vl_logic;
        o_ctrl_trap     : out    vl_logic;
        i_ctrl_misalign : in     vl_logic;
        i_sh_done       : in     vl_logic;
        o_mem_bytecnt   : out    vl_logic_vector(1 downto 0);
        i_mem_misalign  : in     vl_logic;
        i_bne_or_bge    : in     vl_logic;
        i_cond_branch   : in     vl_logic;
        i_dbus_en       : in     vl_logic;
        i_two_stage_op  : in     vl_logic;
        i_branch_op     : in     vl_logic;
        i_shift_op      : in     vl_logic;
        i_sh_right      : in     vl_logic;
        i_alu_rd_sel1   : in     vl_logic;
        i_rd_alu_en     : in     vl_logic;
        i_e_op          : in     vl_logic;
        i_rd_op         : in     vl_logic;
        i_mdu_op        : in     vl_logic;
        o_mdu_valid     : out    vl_logic;
        i_mdu_ready     : in     vl_logic;
        o_dbus_cyc      : out    vl_logic;
        i_dbus_ack      : in     vl_logic;
        o_ibus_cyc      : out    vl_logic;
        i_ibus_ack      : in     vl_logic;
        o_rf_rreq       : out    vl_logic;
        o_rf_wreq       : out    vl_logic;
        i_rf_ready      : in     vl_logic;
        o_rf_rd_en      : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of RESET_STRATEGY : constant is 1;
    attribute mti_svvh_generic_type of WITH_CSR : constant is 2;
    attribute mti_svvh_generic_type of ALIGN : constant is 2;
    attribute mti_svvh_generic_type of MDU : constant is 2;
    attribute mti_svvh_generic_type of W : constant is 1;
end serv_state;
