library verilog;
use verilog.vl_types.all;
entity serv_decode is
    generic(
        PRE_REGISTER    : vl_logic_vector(0 downto 0) := (others => Hi1);
        MDU             : vl_logic_vector(0 downto 0) := (others => Hi0)
    );
    port(
        clk             : in     vl_logic;
        i_wb_rdt        : in     vl_logic_vector(31 downto 2);
        i_wb_en         : in     vl_logic;
        o_sh_right      : out    vl_logic;
        o_bne_or_bge    : out    vl_logic;
        o_cond_branch   : out    vl_logic;
        o_e_op          : out    vl_logic;
        o_ebreak        : out    vl_logic;
        o_branch_op     : out    vl_logic;
        o_shift_op      : out    vl_logic;
        o_rd_op         : out    vl_logic;
        o_two_stage_op  : out    vl_logic;
        o_dbus_en       : out    vl_logic;
        o_mdu_op        : out    vl_logic;
        o_ext_funct3    : out    vl_logic_vector(2 downto 0);
        o_bufreg_rs1_en : out    vl_logic;
        o_bufreg_imm_en : out    vl_logic;
        o_bufreg_clr_lsb: out    vl_logic;
        o_bufreg_sh_signed: out    vl_logic;
        o_ctrl_jal_or_jalr: out    vl_logic;
        o_ctrl_utype    : out    vl_logic;
        o_ctrl_pc_rel   : out    vl_logic;
        o_ctrl_mret     : out    vl_logic;
        o_alu_sub       : out    vl_logic;
        o_alu_bool_op   : out    vl_logic_vector(1 downto 0);
        o_alu_cmp_eq    : out    vl_logic;
        o_alu_cmp_sig   : out    vl_logic;
        o_alu_rd_sel    : out    vl_logic_vector(2 downto 0);
        o_mem_signed    : out    vl_logic;
        o_mem_word      : out    vl_logic;
        o_mem_half      : out    vl_logic;
        o_mem_cmd       : out    vl_logic;
        o_csr_en        : out    vl_logic;
        o_csr_addr      : out    vl_logic_vector(1 downto 0);
        o_csr_mstatus_en: out    vl_logic;
        o_csr_mie_en    : out    vl_logic;
        o_csr_mcause_en : out    vl_logic;
        o_csr_source    : out    vl_logic_vector(1 downto 0);
        o_csr_d_sel     : out    vl_logic;
        o_csr_imm_en    : out    vl_logic;
        o_mtval_pc      : out    vl_logic;
        o_immdec_ctrl   : out    vl_logic_vector(3 downto 0);
        o_immdec_en     : out    vl_logic_vector(3 downto 0);
        o_op_b_source   : out    vl_logic;
        o_rd_mem_en     : out    vl_logic;
        o_rd_csr_en     : out    vl_logic;
        o_rd_alu_en     : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PRE_REGISTER : constant is 2;
    attribute mti_svvh_generic_type of MDU : constant is 2;
end serv_decode;
