library verilog;
use verilog.vl_types.all;
entity serv_top is
    generic(
        WITH_CSR        : integer := 1;
        W               : integer := 1;
        B               : vl_notype;
        PRE_REGISTER    : integer := 1;
        RESET_STRATEGY  : string  := "MINI";
        RESET_PC        : integer := 0;
        DEBUG           : vl_logic_vector(0 downto 0) := (others => Hi0);
        MDU             : vl_logic_vector(0 downto 0) := (others => Hi0);
        COMPRESSED      : vl_logic_vector(0 downto 0) := (others => Hi0);
        ALIGN           : vl_logic_vector(0 downto 0)
    );
    port(
        clk             : in     vl_logic;
        i_rst           : in     vl_logic;
        i_timer_irq     : in     vl_logic;
        o_rf_rreq       : out    vl_logic;
        o_rf_wreq       : out    vl_logic;
        i_rf_ready      : in     vl_logic;
        o_wreg0         : out    vl_logic_vector;
        o_wreg1         : out    vl_logic_vector;
        o_wen0          : out    vl_logic;
        o_wen1          : out    vl_logic;
        o_wdata0        : out    vl_logic_vector;
        o_wdata1        : out    vl_logic_vector;
        o_rreg0         : out    vl_logic_vector;
        o_rreg1         : out    vl_logic_vector;
        i_rdata0        : in     vl_logic_vector;
        i_rdata1        : in     vl_logic_vector;
        o_ibus_adr      : out    vl_logic_vector(31 downto 0);
        o_ibus_cyc      : out    vl_logic;
        i_ibus_rdt      : in     vl_logic_vector(31 downto 0);
        i_ibus_ack      : in     vl_logic;
        o_dbus_adr      : out    vl_logic_vector(31 downto 0);
        o_dbus_dat      : out    vl_logic_vector(31 downto 0);
        o_dbus_sel      : out    vl_logic_vector(3 downto 0);
        o_dbus_we       : out    vl_logic;
        o_dbus_cyc      : out    vl_logic;
        i_dbus_rdt      : in     vl_logic_vector(31 downto 0);
        i_dbus_ack      : in     vl_logic;
        o_ext_funct3    : out    vl_logic_vector(2 downto 0);
        i_ext_ready     : in     vl_logic;
        i_ext_rd        : in     vl_logic_vector(31 downto 0);
        o_ext_rs1       : out    vl_logic_vector(31 downto 0);
        o_ext_rs2       : out    vl_logic_vector(31 downto 0);
        o_mdu_valid     : out    vl_logic;
        o_cnt_done      : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of WITH_CSR : constant is 1;
    attribute mti_svvh_generic_type of W : constant is 1;
    attribute mti_svvh_generic_type of B : constant is 3;
    attribute mti_svvh_generic_type of PRE_REGISTER : constant is 1;
    attribute mti_svvh_generic_type of RESET_STRATEGY : constant is 1;
    attribute mti_svvh_generic_type of RESET_PC : constant is 1;
    attribute mti_svvh_generic_type of DEBUG : constant is 2;
    attribute mti_svvh_generic_type of MDU : constant is 2;
    attribute mti_svvh_generic_type of COMPRESSED : constant is 2;
    attribute mti_svvh_generic_type of ALIGN : constant is 4;
end serv_top;
