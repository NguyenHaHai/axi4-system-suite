library verilog;
use verilog.vl_types.all;
entity serv_axi_wrapper is
    generic(
        ADDR_WIDTH      : integer := 32;
        DATA_WIDTH      : integer := 32;
        ID_WIDTH        : integer := 4;
        WITH_CSR        : integer := 1;
        W               : integer := 1;
        B               : vl_notype;
        PRE_REGISTER    : integer := 1;
        RESET_STRATEGY  : string  := "MINI";
        RESET_PC        : integer := 0;
        DEBUG           : vl_logic_vector(0 downto 0) := (others => Hi0);
        MDU             : vl_logic_vector(0 downto 0) := (others => Hi0);
        COMPRESSED      : vl_logic_vector(0 downto 0) := (others => Hi0);
        ALIGN           : vl_logic_vector(0 downto 0)
    );
    port(
        ACLK            : in     vl_logic;
        ARESETN         : in     vl_logic;
        i_timer_irq     : in     vl_logic;
        M0_AXI_arid     : out    vl_logic_vector;
        M0_AXI_araddr   : out    vl_logic_vector;
        M0_AXI_arlen    : out    vl_logic_vector(7 downto 0);
        M0_AXI_arsize   : out    vl_logic_vector(2 downto 0);
        M0_AXI_arburst  : out    vl_logic_vector(1 downto 0);
        M0_AXI_arlock   : out    vl_logic_vector(1 downto 0);
        M0_AXI_arcache  : out    vl_logic_vector(3 downto 0);
        M0_AXI_arprot   : out    vl_logic_vector(2 downto 0);
        M0_AXI_arqos    : out    vl_logic_vector(3 downto 0);
        M0_AXI_arregion : out    vl_logic_vector(3 downto 0);
        M0_AXI_arvalid  : out    vl_logic;
        M0_AXI_arready  : in     vl_logic;
        M0_AXI_rid      : in     vl_logic_vector;
        M0_AXI_rdata    : in     vl_logic_vector;
        M0_AXI_rresp    : in     vl_logic_vector(1 downto 0);
        M0_AXI_rlast    : in     vl_logic;
        M0_AXI_rvalid   : in     vl_logic;
        M0_AXI_rready   : out    vl_logic;
        M1_AXI_awid     : out    vl_logic_vector;
        M1_AXI_awaddr   : out    vl_logic_vector;
        M1_AXI_awlen    : out    vl_logic_vector(7 downto 0);
        M1_AXI_awsize   : out    vl_logic_vector(2 downto 0);
        M1_AXI_awburst  : out    vl_logic_vector(1 downto 0);
        M1_AXI_awlock   : out    vl_logic_vector(1 downto 0);
        M1_AXI_awcache  : out    vl_logic_vector(3 downto 0);
        M1_AXI_awprot   : out    vl_logic_vector(2 downto 0);
        M1_AXI_awqos    : out    vl_logic_vector(3 downto 0);
        M1_AXI_awregion : out    vl_logic_vector(3 downto 0);
        M1_AXI_awvalid  : out    vl_logic;
        M1_AXI_awready  : in     vl_logic;
        M1_AXI_wdata    : out    vl_logic_vector;
        M1_AXI_wstrb    : out    vl_logic_vector;
        M1_AXI_wlast    : out    vl_logic;
        M1_AXI_wvalid   : out    vl_logic;
        M1_AXI_wready   : in     vl_logic;
        M1_AXI_bid      : in     vl_logic_vector;
        M1_AXI_bresp    : in     vl_logic_vector(1 downto 0);
        M1_AXI_bvalid   : in     vl_logic;
        M1_AXI_bready   : out    vl_logic;
        M1_AXI_arid     : out    vl_logic_vector;
        M1_AXI_araddr   : out    vl_logic_vector;
        M1_AXI_arlen    : out    vl_logic_vector(7 downto 0);
        M1_AXI_arsize   : out    vl_logic_vector(2 downto 0);
        M1_AXI_arburst  : out    vl_logic_vector(1 downto 0);
        M1_AXI_arlock   : out    vl_logic_vector(1 downto 0);
        M1_AXI_arcache  : out    vl_logic_vector(3 downto 0);
        M1_AXI_arprot   : out    vl_logic_vector(2 downto 0);
        M1_AXI_arqos    : out    vl_logic_vector(3 downto 0);
        M1_AXI_arregion : out    vl_logic_vector(3 downto 0);
        M1_AXI_arvalid  : out    vl_logic;
        M1_AXI_arready  : in     vl_logic;
        M1_AXI_rid      : in     vl_logic_vector;
        M1_AXI_rdata    : in     vl_logic_vector;
        M1_AXI_rresp    : in     vl_logic_vector(1 downto 0);
        M1_AXI_rlast    : in     vl_logic;
        M1_AXI_rvalid   : in     vl_logic;
        M1_AXI_rready   : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of WITH_CSR : constant is 1;
    attribute mti_svvh_generic_type of W : constant is 1;
    attribute mti_svvh_generic_type of B : constant is 3;
    attribute mti_svvh_generic_type of PRE_REGISTER : constant is 1;
    attribute mti_svvh_generic_type of RESET_STRATEGY : constant is 1;
    attribute mti_svvh_generic_type of RESET_PC : constant is 1;
    attribute mti_svvh_generic_type of DEBUG : constant is 2;
    attribute mti_svvh_generic_type of MDU : constant is 2;
    attribute mti_svvh_generic_type of COMPRESSED : constant is 2;
    attribute mti_svvh_generic_type of ALIGN : constant is 4;
end serv_axi_wrapper;
