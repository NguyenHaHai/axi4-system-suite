library verilog;
use verilog.vl_types.all;
entity serv_axi_system is
    generic(
        ADDR_WIDTH      : integer := 32;
        DATA_WIDTH      : integer := 32;
        ID_WIDTH        : integer := 4;
        WITH_CSR        : integer := 1;
        W               : integer := 1;
        PRE_REGISTER    : integer := 1;
        RESET_STRATEGY  : string  := "MINI";
        RESET_PC        : integer := 0;
        DEBUG           : vl_logic_vector(0 downto 0) := (others => Hi0);
        MDU             : vl_logic_vector(0 downto 0) := (others => Hi0);
        COMPRESSED      : vl_logic_vector(0 downto 0) := (others => Hi0);
        Num_Of_Slaves   : integer := 2;
        S00_Aw_len      : integer := 8;
        S00_Write_data_bus_width: integer := 32;
        S00_AR_len      : integer := 8;
        S00_Read_data_bus_width: integer := 32;
        S01_Aw_len      : integer := 8;
        S01_Write_data_bus_width: integer := 32;
        S01_AR_len      : integer := 8;
        M00_Aw_len      : integer := 8;
        M00_Write_data_bus_width: integer := 32;
        M00_AR_len      : integer := 8;
        M00_Read_data_bus_width: integer := 32;
        M01_Aw_len      : integer := 8;
        M01_AR_len      : integer := 8;
        Is_Master_AXI_4 : vl_logic := Hi1;
        Num_Of_Masters  : integer := 2;
        Master_ID_Width : integer := 1;
        AXI4_AR_len     : integer := 8;
        SLAVE0_ADDR1    : integer := 0;
        SLAVE0_ADDR2    : integer := 1073741823;
        SLAVE1_ADDR1    : integer := 1073741824;
        SLAVE1_ADDR2    : integer := 2147483647
    );
    port(
        ACLK            : in     vl_logic;
        ARESETN         : in     vl_logic;
        i_timer_irq     : in     vl_logic;
        M00_AXI_araddr  : out    vl_logic_vector;
        M00_AXI_arlen   : out    vl_logic_vector(7 downto 0);
        M00_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M00_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M00_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M00_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M00_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M00_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M00_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M00_AXI_arvalid : out    vl_logic;
        M00_AXI_arready : in     vl_logic;
        M00_AXI_rdata   : in     vl_logic_vector;
        M00_AXI_rresp   : in     vl_logic_vector(1 downto 0);
        M00_AXI_rlast   : in     vl_logic;
        M00_AXI_rvalid  : in     vl_logic;
        M00_AXI_rready  : out    vl_logic;
        M01_AXI_awid    : out    vl_logic_vector;
        M01_AXI_awaddr  : out    vl_logic_vector;
        M01_AXI_awlen   : out    vl_logic_vector(7 downto 0);
        M01_AXI_awsize  : out    vl_logic_vector(2 downto 0);
        M01_AXI_awburst : out    vl_logic_vector(1 downto 0);
        M01_AXI_awlock  : out    vl_logic_vector(1 downto 0);
        M01_AXI_awcache : out    vl_logic_vector(3 downto 0);
        M01_AXI_awprot  : out    vl_logic_vector(2 downto 0);
        M01_AXI_awqos   : out    vl_logic_vector(3 downto 0);
        M01_AXI_awregion: out    vl_logic_vector(3 downto 0);
        M01_AXI_awvalid : out    vl_logic;
        M01_AXI_awready : in     vl_logic;
        M01_AXI_wdata   : out    vl_logic_vector;
        M01_AXI_wstrb   : out    vl_logic_vector;
        M01_AXI_wlast   : out    vl_logic;
        M01_AXI_wvalid  : out    vl_logic;
        M01_AXI_wready  : in     vl_logic;
        M01_AXI_bid     : in     vl_logic_vector;
        M01_AXI_bresp   : in     vl_logic_vector(1 downto 0);
        M01_AXI_bvalid  : in     vl_logic;
        M01_AXI_bready  : out    vl_logic;
        M01_AXI_arid    : out    vl_logic_vector;
        M01_AXI_araddr  : out    vl_logic_vector;
        M01_AXI_arlen   : out    vl_logic_vector(7 downto 0);
        M01_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M01_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M01_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M01_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M01_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M01_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M01_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M01_AXI_arvalid : out    vl_logic;
        M01_AXI_arready : in     vl_logic;
        M01_AXI_rid     : in     vl_logic_vector;
        M01_AXI_rdata   : in     vl_logic_vector;
        M01_AXI_rresp   : in     vl_logic_vector(1 downto 0);
        M01_AXI_rlast   : in     vl_logic;
        M01_AXI_rvalid  : in     vl_logic;
        M01_AXI_rready  : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of WITH_CSR : constant is 1;
    attribute mti_svvh_generic_type of W : constant is 1;
    attribute mti_svvh_generic_type of PRE_REGISTER : constant is 1;
    attribute mti_svvh_generic_type of RESET_STRATEGY : constant is 1;
    attribute mti_svvh_generic_type of RESET_PC : constant is 1;
    attribute mti_svvh_generic_type of DEBUG : constant is 2;
    attribute mti_svvh_generic_type of MDU : constant is 2;
    attribute mti_svvh_generic_type of COMPRESSED : constant is 2;
    attribute mti_svvh_generic_type of Num_Of_Slaves : constant is 1;
    attribute mti_svvh_generic_type of S00_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of S00_Write_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of S00_AR_len : constant is 1;
    attribute mti_svvh_generic_type of S00_Read_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of S01_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of S01_Write_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of S01_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M00_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M00_Write_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of M00_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M00_Read_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of M01_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M01_AR_len : constant is 1;
    attribute mti_svvh_generic_type of Is_Master_AXI_4 : constant is 1;
    attribute mti_svvh_generic_type of Num_Of_Masters : constant is 1;
    attribute mti_svvh_generic_type of Master_ID_Width : constant is 1;
    attribute mti_svvh_generic_type of AXI4_AR_len : constant is 1;
    attribute mti_svvh_generic_type of SLAVE0_ADDR1 : constant is 1;
    attribute mti_svvh_generic_type of SLAVE0_ADDR2 : constant is 1;
    attribute mti_svvh_generic_type of SLAVE1_ADDR1 : constant is 1;
    attribute mti_svvh_generic_type of SLAVE1_ADDR2 : constant is 1;
end serv_axi_system;
