library verilog;
use verilog.vl_types.all;
entity AXI_Interconnect_2S_RDONLY is
    port(
        ACLK            : in     vl_logic;
        ARESETN         : in     vl_logic;
        S00_AXI_araddr  : in     vl_logic_vector(31 downto 0);
        S00_AXI_arlen   : in     vl_logic_vector(7 downto 0);
        S00_AXI_arsize  : in     vl_logic_vector(2 downto 0);
        S00_AXI_arburst : in     vl_logic_vector(1 downto 0);
        S00_AXI_arlock  : in     vl_logic_vector(1 downto 0);
        S00_AXI_arcache : in     vl_logic_vector(3 downto 0);
        S00_AXI_arprot  : in     vl_logic_vector(2 downto 0);
        S00_AXI_arregion: in     vl_logic_vector(3 downto 0);
        S00_AXI_arqos   : in     vl_logic_vector(3 downto 0);
        S00_AXI_arvalid : in     vl_logic;
        S00_AXI_arready : out    vl_logic;
        S00_AXI_rdata   : out    vl_logic_vector(31 downto 0);
        S00_AXI_rresp   : out    vl_logic_vector(1 downto 0);
        S00_AXI_rlast   : out    vl_logic;
        S00_AXI_rvalid  : out    vl_logic;
        S00_AXI_rready  : in     vl_logic;
        S01_AXI_araddr  : in     vl_logic_vector(31 downto 0);
        S01_AXI_arlen   : in     vl_logic_vector(7 downto 0);
        S01_AXI_arsize  : in     vl_logic_vector(2 downto 0);
        S01_AXI_arburst : in     vl_logic_vector(1 downto 0);
        S01_AXI_arlock  : in     vl_logic_vector(1 downto 0);
        S01_AXI_arcache : in     vl_logic_vector(3 downto 0);
        S01_AXI_arprot  : in     vl_logic_vector(2 downto 0);
        S01_AXI_arregion: in     vl_logic_vector(3 downto 0);
        S01_AXI_arqos   : in     vl_logic_vector(3 downto 0);
        S01_AXI_arvalid : in     vl_logic;
        S01_AXI_arready : out    vl_logic;
        S01_AXI_rdata   : out    vl_logic_vector(31 downto 0);
        S01_AXI_rresp   : out    vl_logic_vector(1 downto 0);
        S01_AXI_rlast   : out    vl_logic;
        S01_AXI_rvalid  : out    vl_logic;
        S01_AXI_rready  : in     vl_logic;
        M00_AXI_araddr  : out    vl_logic_vector(31 downto 0);
        M00_AXI_arlen   : out    vl_logic_vector(7 downto 0);
        M00_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M00_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M00_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M00_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M00_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M00_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M00_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M00_AXI_arvalid : out    vl_logic;
        M00_AXI_arready : in     vl_logic;
        M00_AXI_rdata   : in     vl_logic_vector(31 downto 0);
        M00_AXI_rresp   : in     vl_logic_vector(1 downto 0);
        M00_AXI_rlast   : in     vl_logic;
        M00_AXI_rvalid  : in     vl_logic;
        M00_AXI_rready  : out    vl_logic;
        M01_AXI_araddr  : out    vl_logic_vector(31 downto 0);
        M01_AXI_arlen   : out    vl_logic_vector(7 downto 0);
        M01_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M01_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M01_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M01_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M01_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M01_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M01_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M01_AXI_arvalid : out    vl_logic;
        M01_AXI_arready : in     vl_logic;
        M01_AXI_rdata   : in     vl_logic_vector(31 downto 0);
        M01_AXI_rresp   : in     vl_logic_vector(1 downto 0);
        M01_AXI_rlast   : in     vl_logic;
        M01_AXI_rvalid  : in     vl_logic;
        M01_AXI_rready  : out    vl_logic;
        slave0_addr1    : in     vl_logic_vector(31 downto 0);
        slave0_addr2    : in     vl_logic_vector(31 downto 0);
        slave1_addr1    : in     vl_logic_vector(31 downto 0);
        slave1_addr2    : in     vl_logic_vector(31 downto 0)
    );
end AXI_Interconnect_2S_RDONLY;
